//-----------------------------------------------------------------
//                      FPGA Media Player
//                            V0.1
//                     Ultra-Embedded.com
//                        Copyright 2020
//
//                   admin@ultra-embedded.com
//
//                     License: Apache 2.0
//-----------------------------------------------------------------
// Copyright 2020 Ultra-Embedded.com
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//-----------------------------------------------------------------

module bootrom
(
    // Inputs
     input           clk_i
    ,input           rst_i
    ,input           inport_awvalid_i
    ,input  [ 31:0]  inport_awaddr_i
    ,input  [  3:0]  inport_awid_i
    ,input  [  7:0]  inport_awlen_i
    ,input  [  1:0]  inport_awburst_i
    ,input           inport_wvalid_i
    ,input  [ 31:0]  inport_wdata_i
    ,input  [  3:0]  inport_wstrb_i
    ,input           inport_wlast_i
    ,input           inport_bready_i
    ,input           inport_arvalid_i
    ,input  [ 31:0]  inport_araddr_i
    ,input  [  3:0]  inport_arid_i
    ,input  [  7:0]  inport_arlen_i
    ,input  [  1:0]  inport_arburst_i
    ,input           inport_rready_i

    // Outputs
    ,output          inport_awready_o
    ,output          inport_wready_o
    ,output          inport_bvalid_o
    ,output [  1:0]  inport_bresp_o
    ,output [  3:0]  inport_bid_o
    ,output          inport_arready_o
    ,output          inport_rvalid_o
    ,output [ 31:0]  inport_rdata_o
    ,output [  1:0]  inport_rresp_o
    ,output [  3:0]  inport_rid_o
    ,output          inport_rlast_o
);



//-----------------------------------------------------------------
// AXI logic
//-----------------------------------------------------------------
wire [  3:0]  ram_wr_w;
wire          ram_rd_w;
wire [ 31:0]  ram_addr_w;
wire [ 31:0]  ram_write_data_w;
wire [ 31:0]  ram_read_data_w;

bootrom_bridge
u_axi
(
    // Inputs
    .clk_i(clk_i),
    .rst_i(rst_i),
    .axi_awvalid_i(inport_awvalid_i),
    .axi_awaddr_i(inport_awaddr_i),
    .axi_awid_i(inport_awid_i),
    .axi_awlen_i(inport_awlen_i),
    .axi_awburst_i(inport_awburst_i),
    .axi_wvalid_i(inport_wvalid_i),
    .axi_wdata_i(inport_wdata_i),
    .axi_wstrb_i(inport_wstrb_i),
    .axi_wlast_i(inport_wlast_i),
    .axi_bready_i(inport_bready_i),
    .axi_arvalid_i(inport_arvalid_i),
    .axi_araddr_i(inport_araddr_i),
    .axi_arid_i(inport_arid_i),
    .axi_arlen_i(inport_arlen_i),
    .axi_arburst_i(inport_arburst_i),
    .axi_rready_i(inport_rready_i),
    .ram_read_data_i(ram_read_data_w),
    .ram_accept_i(1'b1),

    // Outputs
    .axi_awready_o(inport_awready_o),
    .axi_wready_o(inport_wready_o),
    .axi_bvalid_o(inport_bvalid_o),
    .axi_bresp_o(inport_bresp_o),
    .axi_bid_o(inport_bid_o),
    .axi_arready_o(inport_arready_o),
    .axi_rvalid_o(inport_rvalid_o),
    .axi_rdata_o(inport_rdata_o),
    .axi_rresp_o(inport_rresp_o),
    .axi_rid_o(inport_rid_o),
    .axi_rlast_o(inport_rlast_o),
    .ram_wr_o(ram_wr_w),
    .ram_rd_o(ram_rd_w),
    .ram_addr_o(ram_addr_w),
    .ram_write_data_o(ram_write_data_w)
);

//-----------------------------------------------------------------
// RAM 8KB
//-----------------------------------------------------------------
wire [10:0] addr_w = ram_addr_w[12:2];

reg [31:0] ram [2047:0] /*verilator public*/;

reg [31:0] ram_read_q;

initial
begin
    ram[0] = 32'h980006f;
    ram[1] = 32'h0;
    ram[2] = 32'h0;
    ram[3] = 32'h0;
    ram[4] = 32'h880006f;
    ram[5] = 32'h0;
    ram[6] = 32'h0;
    ram[7] = 32'h0;
    ram[8] = 32'h0;
    ram[9] = 32'h0;
    ram[10] = 32'h0;
    ram[11] = 32'h0;
    ram[12] = 32'h0;
    ram[13] = 32'h0;
    ram[14] = 32'h0;
    ram[15] = 32'h0;
    ram[16] = 32'h0;
    ram[17] = 32'h0;
    ram[18] = 32'hfe010113;
    ram[19] = 32'h1112e23;
    ram[20] = 32'h1012c23;
    ram[21] = 32'hf12a23;
    ram[22] = 32'he12823;
    ram[23] = 32'hd12623;
    ram[24] = 32'hc12423;
    ram[25] = 32'hb12223;
    ram[26] = 32'ha12023;
    ram[27] = 32'h820005b7;
    ram[28] = 32'h1458593;
    ram[29] = 32'h25a223;
    ram[30] = 32'h55a023;
    ram[31] = 32'h3a159073;
    ram[32] = 32'h3a259073;
    ram[33] = 32'h5a283;
    ram[34] = 32'hfe029ce3;
    ram[35] = 32'h12503;
    ram[36] = 32'h2010113;
    ram[37] = 32'h8067;
    ram[38] = 32'h82002137;
    ram[39] = 32'h8e810113;
    ram[40] = 32'h820002b7;
    ram[41] = 32'h2028293;
    ram[42] = 32'h82002337;
    ram[43] = 32'h8f830313;
    ram[44] = 32'h2a023;
    ram[45] = 32'h428293;
    ram[46] = 32'hfe62cce3;
    ram[47] = 32'h820002b7;
    ram[48] = 32'h28293;
    ram[49] = 32'h82000337;
    ram[50] = 32'h2030313;
    ram[51] = 32'h400023b7;
    ram[52] = 32'hefc38393;
    ram[53] = 32'h3ae03;
    ram[54] = 32'h1c2a023;
    ram[55] = 32'h428293;
    ram[56] = 32'h438393;
    ram[57] = 32'hfe62c8e3;
    ram[58] = 32'h4d5010ef;
    ram[59] = 32'h517;
    ram[60] = 32'hf4850513;
    ram[61] = 32'h52503;
    ram[62] = 32'h597;
    ram[63] = 32'hf4058593;
    ram[64] = 32'h28000ef;
    ram[65] = 32'h4000ef;
    ram[66] = 32'hffc10113;
    ram[67] = 32'h112023;
    ram[68] = 32'h297;
    ram[69] = 32'hff828293;
    ram[70] = 32'hf31ff0ef;
    ram[71] = 32'h12083;
    ram[72] = 32'h410113;
    ram[73] = 32'h8067;
    ram[74] = 32'h40002537;
    ram[75] = 32'hff010113;
    ram[76] = 32'he7850513;
    ram[77] = 32'h112623;
    ram[78] = 32'h812423;
    ram[79] = 32'h912223;
    ram[80] = 32'h1212023;
    ram[81] = 32'h485010ef;
    ram[82] = 32'h1dc000ef;
    ram[83] = 32'h2055263;
    ram[84] = 32'hfff00413;
    ram[85] = 32'h40513;
    ram[86] = 32'hc12083;
    ram[87] = 32'h812403;
    ram[88] = 32'h412483;
    ram[89] = 32'h12903;
    ram[90] = 32'h1010113;
    ram[91] = 32'h8067;
    ram[92] = 32'h3fc010ef;
    ram[93] = 32'h40000537;
    ram[94] = 32'h593;
    ram[95] = 32'h55850513;
    ram[96] = 32'h43c010ef;
    ram[97] = 32'h50413;
    ram[98] = 32'hfc0514e3;
    ram[99] = 32'h400025b7;
    ram[100] = 32'h40002537;
    ram[101] = 32'he8858593;
    ram[102] = 32'he8c50513;
    ram[103] = 32'h47c010ef;
    ram[104] = 32'h50493;
    ram[105] = 32'hfa0506e3;
    ram[106] = 32'h80000937;
    ram[107] = 32'h48693;
    ram[108] = 32'h8637;
    ram[109] = 32'h100593;
    ram[110] = 32'h90513;
    ram[111] = 32'h674010ef;
    ram[112] = 32'ha05663;
    ram[113] = 32'ha90933;
    ram[114] = 32'hfe5ff06f;
    ram[115] = 32'h48513;
    ram[116] = 32'h5b8010ef;
    ram[117] = 32'h3a001073;
    ram[118] = 32'h100f;
    ram[119] = 32'h13;
    ram[120] = 32'h13;
    ram[121] = 32'h13;
    ram[122] = 32'h800007b7;
    ram[123] = 32'h780e7;
    ram[124] = 32'hf65ff06f;
    ram[125] = 32'h185d713;
    ram[126] = 32'h47b7;
    ram[127] = 32'he7e7b3;
    ram[128] = 32'h851713;
    ram[129] = 32'h859593;
    ram[130] = 32'he7e7b3;
    ram[131] = 32'hfe010113;
    ram[132] = 32'h1079793;
    ram[133] = 32'h105d713;
    ram[134] = 32'h912a23;
    ram[135] = 32'h112e23;
    ram[136] = 32'h812c23;
    ram[137] = 32'h1212823;
    ram[138] = 32'h1312623;
    ram[139] = 32'he7e733;
    ram[140] = 32'h960007b7;
    ram[141] = 32'he7a623;
    ram[142] = 32'hb7a823;
    ram[143] = 32'h60493;
    ram[144] = 32'h800007b7;
    ram[145] = 32'h8061063;
    ram[146] = 32'hfef50713;
    ram[147] = 32'h100693;
    ram[148] = 32'hce6e063;
    ram[149] = 32'h47e793;
    ram[150] = 32'h82001737;
    ram[151] = 32'h8d072703;
    ram[152] = 32'h70463;
    ram[153] = 32'h87e793;
    ram[154] = 32'h1200713;
    ram[155] = 32'h6e51063;
    ram[156] = 32'h8737;
    ram[157] = 32'hf0070713;
    ram[158] = 32'he7e7b3;
    ram[159] = 32'h96000737;
    ram[160] = 32'hf72023;
    ram[161] = 32'h3ad010ef;
    ram[162] = 32'h50913;
    ram[163] = 32'h96000437;
    ram[164] = 32'hfa00993;
    ram[165] = 32'h842783;
    ram[166] = 32'h17f793;
    ram[167] = 32'h4079063;
    ram[168] = 32'h100513;
    ram[169] = 32'h4048863;
    ram[170] = 32'h1442783;
    ram[171] = 32'h87d713;
    ram[172] = 32'h1842783;
    ram[173] = 32'h1879793;
    ram[174] = 32'he7e7b3;
    ram[175] = 32'hf4a023;
    ram[176] = 32'h340006f;
    ram[177] = 32'h178793;
    ram[178] = 32'hf81ff06f;
    ram[179] = 32'h1800713;
    ram[180] = 32'hfae516e3;
    ram[181] = 32'h207e793;
    ram[182] = 32'hfa5ff06f;
    ram[183] = 32'h355010ef;
    ram[184] = 32'h41250533;
    ram[185] = 32'hfaa9d8e3;
    ram[186] = 32'h400007b7;
    ram[187] = 32'hf42023;
    ram[188] = 32'h513;
    ram[189] = 32'h1c12083;
    ram[190] = 32'h1812403;
    ram[191] = 32'h1412483;
    ram[192] = 32'h1012903;
    ram[193] = 32'hc12983;
    ram[194] = 32'h2010113;
    ram[195] = 32'h8067;
    ram[196] = 32'h1800713;
    ram[197] = 32'hf4e502e3;
    ram[198] = 32'h1200713;
    ram[199] = 32'hf6e510e3;
    ram[200] = 32'hf51ff06f;
    ram[201] = 32'hfe010113;
    ram[202] = 32'h812c23;
    ram[203] = 32'h912a23;
    ram[204] = 32'h112e23;
    ram[205] = 32'h1212823;
    ram[206] = 32'h960007b7;
    ram[207] = 32'h100713;
    ram[208] = 32'he7a223;
    ram[209] = 32'h613;
    ram[210] = 32'h593;
    ram[211] = 32'h513;
    ram[212] = 32'hea5ff0ef;
    ram[213] = 32'h413;
    ram[214] = 32'h400493;
    ram[215] = 32'hc10613;
    ram[216] = 32'h1aa00593;
    ram[217] = 32'h800513;
    ram[218] = 32'he8dff0ef;
    ram[219] = 32'h51863;
    ram[220] = 32'h140793;
    ram[221] = 32'h84ca63;
    ram[222] = 32'h78413;
    ram[223] = 32'hc12703;
    ram[224] = 32'h1aa00793;
    ram[225] = 32'hfcf71ce3;
    ram[226] = 32'h82001437;
    ram[227] = 32'hc10613;
    ram[228] = 32'h593;
    ram[229] = 32'h3700513;
    ram[230] = 32'he5dff0ef;
    ram[231] = 32'hc10613;
    ram[232] = 32'h401005b7;
    ram[233] = 32'h2900513;
    ram[234] = 32'he4dff0ef;
    ram[235] = 32'hc12703;
    ram[236] = 32'h1e75793;
    ram[237] = 32'h17f793;
    ram[238] = 32'h8cf42623;
    ram[239] = 32'hfc0758e3;
    ram[240] = 32'h960007b7;
    ram[241] = 32'h42000737;
    ram[242] = 32'he7a623;
    ram[243] = 32'h80000737;
    ram[244] = 32'h7a823;
    ram[245] = 32'h270713;
    ram[246] = 32'he7a023;
    ram[247] = 32'h255010ef;
    ram[248] = 32'h50493;
    ram[249] = 32'h96000437;
    ram[250] = 32'hfa00913;
    ram[251] = 32'h842783;
    ram[252] = 32'h17f793;
    ram[253] = 32'h79e63;
    ram[254] = 32'h1442783;
    ram[255] = 32'h1842783;
    ram[256] = 32'h1c42783;
    ram[257] = 32'h2042783;
    ram[258] = 32'h2442783;
    ram[259] = 32'h180006f;
    ram[260] = 32'h221010ef;
    ram[261] = 32'h40950533;
    ram[262] = 32'hfca95ae3;
    ram[263] = 32'h400007b7;
    ram[264] = 32'hf42023;
    ram[265] = 32'hc10613;
    ram[266] = 32'h593;
    ram[267] = 32'h300513;
    ram[268] = 32'hdc5ff0ef;
    ram[269] = 32'hc12783;
    ram[270] = 32'hffff0437;
    ram[271] = 32'hc10613;
    ram[272] = 32'hf47433;
    ram[273] = 32'h40593;
    ram[274] = 32'hd00513;
    ram[275] = 32'hda9ff0ef;
    ram[276] = 32'hc12783;
    ram[277] = 32'h2737;
    ram[278] = 32'he0070713;
    ram[279] = 32'he7f7b3;
    ram[280] = 32'h80078713;
    ram[281] = 32'h6070063;
    ram[282] = 32'h1737;
    ram[283] = 32'h80070693;
    ram[284] = 32'h4f6e063;
    ram[285] = 32'h20000713;
    ram[286] = 32'hae78e63;
    ram[287] = 32'hf76863;
    ram[288] = 32'ha078a63;
    ram[289] = 32'h20100693;
    ram[290] = 32'hb00006f;
    ram[291] = 32'h40000713;
    ram[292] = 32'hae78263;
    ram[293] = 32'h60000713;
    ram[294] = 32'hfee796e3;
    ram[295] = 32'hc10613;
    ram[296] = 32'h40593;
    ram[297] = 32'h700513;
    ram[298] = 32'hd4dff0ef;
    ram[299] = 32'h180006f;
    ram[300] = 32'hc0070693;
    ram[301] = 32'hd78863;
    ram[302] = 32'h6f6e463;
    ram[303] = 32'ha0070713;
    ram[304] = 32'hfce792e3;
    ram[305] = 32'h6400513;
    ram[306] = 32'h145010ef;
    ram[307] = 32'hc10613;
    ram[308] = 32'h40593;
    ram[309] = 32'h3700513;
    ram[310] = 32'hd1dff0ef;
    ram[311] = 32'hc10613;
    ram[312] = 32'h200593;
    ram[313] = 32'h600513;
    ram[314] = 32'hd0dff0ef;
    ram[315] = 32'h40002537;
    ram[316] = 32'h820017b7;
    ram[317] = 32'h100713;
    ram[318] = 32'hecc50513;
    ram[319] = 32'h8ce7a823;
    ram[320] = 32'h61010ef;
    ram[321] = 32'h1c12083;
    ram[322] = 32'h1812403;
    ram[323] = 32'h1412483;
    ram[324] = 32'h1012903;
    ram[325] = 32'h100513;
    ram[326] = 32'h2010113;
    ram[327] = 32'h8067;
    ram[328] = 32'he0070693;
    ram[329] = 32'hd78463;
    ram[330] = 32'hf4e79ee3;
    ram[331] = 32'h1fd00693;
    ram[332] = 32'h80006f;
    ram[333] = 32'h1e900693;
    ram[334] = 32'h40002637;
    ram[335] = 32'h400025b7;
    ram[336] = 32'h40002537;
    ram[337] = 32'he9860613;
    ram[338] = 32'heb458593;
    ram[339] = 32'hec450513;
    ram[340] = 32'had010ef;
    ram[341] = 32'hf71ff06f;
    ram[342] = 32'h18060463;
    ram[343] = 32'hfb010113;
    ram[344] = 32'h3412c23;
    ram[345] = 32'h3512a23;
    ram[346] = 32'h951a13;
    ram[347] = 32'h5ab7;
    ram[348] = 32'h4812423;
    ram[349] = 32'h4912223;
    ram[350] = 32'h5212023;
    ram[351] = 32'h3312e23;
    ram[352] = 32'h3612823;
    ram[353] = 32'h3712623;
    ram[354] = 32'h3812423;
    ram[355] = 32'h3912223;
    ram[356] = 32'h3a12023;
    ram[357] = 32'h4112623;
    ram[358] = 32'h1b12e23;
    ram[359] = 32'h50493;
    ram[360] = 32'h58913;
    ram[361] = 32'ha609b3;
    ram[362] = 32'h40ba0a33;
    ram[363] = 32'h82001b37;
    ram[364] = 32'h40002bb7;
    ram[365] = 32'h40002c37;
    ram[366] = 32'h40002cb7;
    ram[367] = 32'h100a8a93;
    ram[368] = 32'h96000437;
    ram[369] = 32'h82001d37;
    ram[370] = 32'h5349263;
    ram[371] = 32'h4c12083;
    ram[372] = 32'h4812403;
    ram[373] = 32'h4412483;
    ram[374] = 32'h4012903;
    ram[375] = 32'h3c12983;
    ram[376] = 32'h3812a03;
    ram[377] = 32'h3412a83;
    ram[378] = 32'h3012b03;
    ram[379] = 32'h2c12b83;
    ram[380] = 32'h2812c03;
    ram[381] = 32'h2412c83;
    ram[382] = 32'h2012d03;
    ram[383] = 32'h1c12d83;
    ram[384] = 32'h100513;
    ram[385] = 32'h5010113;
    ram[386] = 32'h8067;
    ram[387] = 32'h8ccb2783;
    ram[388] = 32'h48d93;
    ram[389] = 32'h79463;
    ram[390] = 32'h1490db3;
    ram[391] = 32'h397793;
    ram[392] = 32'h78c63;
    ram[393] = 32'h15900693;
    ram[394] = 32'he98b8613;
    ram[395] = 32'hee0c0593;
    ram[396] = 32'hec4c8513;
    ram[397] = 32'h7c8010ef;
    ram[398] = 32'h18dd793;
    ram[399] = 32'h157e7b3;
    ram[400] = 32'h8d9d93;
    ram[401] = 32'h1079793;
    ram[402] = 32'h10dd713;
    ram[403] = 32'he7e733;
    ram[404] = 32'h8d0d2783;
    ram[405] = 32'he42623;
    ram[406] = 32'h1b42823;
    ram[407] = 32'h4078863;
    ram[408] = 32'h800007b7;
    ram[409] = 32'hd78793;
    ram[410] = 32'hf42023;
    ram[411] = 32'h7c4010ef;
    ram[412] = 32'h50d93;
    ram[413] = 32'h3e800713;
    ram[414] = 32'h842783;
    ram[415] = 32'h17f793;
    ram[416] = 32'h2079c63;
    ram[417] = 32'h1442783;
    ram[418] = 32'h1842783;
    ram[419] = 32'h90713;
    ram[420] = 32'h842783;
    ram[421] = 32'h87f793;
    ram[422] = 32'h2079e63;
    ram[423] = 32'h2c42783;
    ram[424] = 32'h470713;
    ram[425] = 32'hfef72e23;
    ram[426] = 32'hfe9ff06f;
    ram[427] = 32'h800007b7;
    ram[428] = 32'h578793;
    ram[429] = 32'hfb5ff06f;
    ram[430] = 32'he12623;
    ram[431] = 32'h774010ef;
    ram[432] = 32'hc12703;
    ram[433] = 32'h41b50533;
    ram[434] = 32'hfaa758e3;
    ram[435] = 32'h400007b7;
    ram[436] = 32'hf42023;
    ram[437] = 32'h20090913;
    ram[438] = 32'h148493;
    ram[439] = 32'heedff06f;
    ram[440] = 32'h100513;
    ram[441] = 32'h8067;
    ram[442] = 32'h100513;
    ram[443] = 32'h8067;
    ram[444] = 32'h513;
    ram[445] = 32'h8067;
    ram[446] = 32'h100513;
    ram[447] = 32'h8067;
    ram[448] = 32'hff010113;
    ram[449] = 32'h812423;
    ram[450] = 32'h112623;
    ram[451] = 32'h912223;
    ram[452] = 32'hfff00793;
    ram[453] = 32'h24f52223;
    ram[454] = 32'h24052423;
    ram[455] = 32'h2052223;
    ram[456] = 32'h50413;
    ram[457] = 32'h42c010ef;
    ram[458] = 32'h3442783;
    ram[459] = 32'h79e63;
    ram[460] = 32'hfff00513;
    ram[461] = 32'hc12083;
    ram[462] = 32'h812403;
    ram[463] = 32'h412483;
    ram[464] = 32'h1010113;
    ram[465] = 32'h8067;
    ram[466] = 32'h4440493;
    ram[467] = 32'h100613;
    ram[468] = 32'h48593;
    ram[469] = 32'h513;
    ram[470] = 32'h780e7;
    ram[471] = 32'hfc050ae3;
    ram[472] = 32'h24042703;
    ram[473] = 32'hffff07b7;
    ram[474] = 32'he7f7b3;
    ram[475] = 32'haa550737;
    ram[476] = 32'he78663;
    ram[477] = 32'hffd00513;
    ram[478] = 32'hfbdff06f;
    ram[479] = 32'h24344783;
    ram[480] = 32'h24244703;
    ram[481] = 32'hffc00513;
    ram[482] = 32'h879793;
    ram[483] = 32'he787b3;
    ram[484] = 32'hb737;
    ram[485] = 32'ha5570713;
    ram[486] = 32'hf8e79ee3;
    ram[487] = 32'h20644703;
    ram[488] = 32'hf00793;
    ram[489] = 32'h22e7ea63;
    ram[490] = 32'h100793;
    ram[491] = 32'he6b7;
    ram[492] = 32'he797b3;
    ram[493] = 32'h86068693;
    ram[494] = 32'hd7f7b3;
    ram[495] = 32'h79863;
    ram[496] = 32'h20070c63;
    ram[497] = 32'h600793;
    ram[498] = 32'h20e7e863;
    ram[499] = 32'h20d44783;
    ram[500] = 32'h20c44703;
    ram[501] = 32'h1879793;
    ram[502] = 32'h1071713;
    ram[503] = 32'he787b3;
    ram[504] = 32'h20a44703;
    ram[505] = 32'he787b3;
    ram[506] = 32'h20b44703;
    ram[507] = 32'h871713;
    ram[508] = 32'he787b3;
    ram[509] = 32'hf42e23;
    ram[510] = 32'h3442783;
    ram[511] = 32'h1c42503;
    ram[512] = 32'h100613;
    ram[513] = 32'h48593;
    ram[514] = 32'h780e7;
    ram[515] = 32'hf20502e3;
    ram[516] = 32'h5044783;
    ram[517] = 32'h4f44703;
    ram[518] = 32'hffe00513;
    ram[519] = 32'h879793;
    ram[520] = 32'he787b3;
    ram[521] = 32'h20000713;
    ram[522] = 32'hf0e796e3;
    ram[523] = 32'h5344583;
    ram[524] = 32'h5244e03;
    ram[525] = 32'h5644603;
    ram[526] = 32'h5544683;
    ram[527] = 32'h859593;
    ram[528] = 32'h1c58533;
    ram[529] = 32'h861613;
    ram[530] = 32'h5b44703;
    ram[531] = 32'h1051e93;
    ram[532] = 32'h5144303;
    ram[533] = 32'hd60533;
    ram[534] = 32'h5a44783;
    ram[535] = 32'h1051513;
    ram[536] = 32'h1055513;
    ram[537] = 32'h871713;
    ram[538] = 32'h640023;
    ram[539] = 32'h2a41423;
    ram[540] = 32'hf70733;
    ram[541] = 32'h10ede93;
    ram[542] = 32'h5444883;
    ram[543] = 32'h16070263;
    ram[544] = 32'h2e42023;
    ram[545] = 32'h7344803;
    ram[546] = 32'h7244783;
    ram[547] = 32'h551513;
    ram[548] = 32'h1881813;
    ram[549] = 32'h1079793;
    ram[550] = 32'hf80833;
    ram[551] = 32'h7044783;
    ram[552] = 32'h1ff50513;
    ram[553] = 32'h40955513;
    ram[554] = 32'hf80833;
    ram[555] = 32'h7144783;
    ram[556] = 32'ha42823;
    ram[557] = 32'h1c42503;
    ram[558] = 32'h879793;
    ram[559] = 32'hf80833;
    ram[560] = 32'h7544783;
    ram[561] = 32'h1042423;
    ram[562] = 32'h7444803;
    ram[563] = 32'h879793;
    ram[564] = 32'hae8533;
    ram[565] = 32'h10787b3;
    ram[566] = 32'hf41c23;
    ram[567] = 32'h2042783;
    ram[568] = 32'ha42a23;
    ram[569] = 32'h2f887b3;
    ram[570] = 32'hfe8833;
    ram[571] = 32'ha787b3;
    ram[572] = 32'hf42223;
    ram[573] = 32'h24344783;
    ram[574] = 32'h24244503;
    ram[575] = 32'h1042623;
    ram[576] = 32'h879793;
    ram[577] = 32'ha787b3;
    ram[578] = 32'hb537;
    ram[579] = 32'ha5550513;
    ram[580] = 32'he6a792e3;
    ram[581] = 32'hd60633;
    ram[582] = 32'h561613;
    ram[583] = 32'h1ff60613;
    ram[584] = 32'h40965613;
    ram[585] = 32'h70693;
    ram[586] = 32'h2071663;
    ram[587] = 32'h6b44683;
    ram[588] = 32'h6a44703;
    ram[589] = 32'h1869693;
    ram[590] = 32'h1071713;
    ram[591] = 32'he686b3;
    ram[592] = 32'h6844703;
    ram[593] = 32'he686b3;
    ram[594] = 32'h6944703;
    ram[595] = 32'h871713;
    ram[596] = 32'he686b3;
    ram[597] = 32'h5844703;
    ram[598] = 32'h5744783;
    ram[599] = 32'h871713;
    ram[600] = 32'hf70733;
    ram[601] = 32'h2071663;
    ram[602] = 32'h6744703;
    ram[603] = 32'h6644783;
    ram[604] = 32'h1871713;
    ram[605] = 32'h1079793;
    ram[606] = 32'hf70733;
    ram[607] = 32'h6444783;
    ram[608] = 32'hf70733;
    ram[609] = 32'h6544783;
    ram[610] = 32'h879793;
    ram[611] = 32'hf70733;
    ram[612] = 32'h2d886b3;
    ram[613] = 32'h1c587b3;
    ram[614] = 32'hc787b3;
    ram[615] = 32'hffb00513;
    ram[616] = 32'hd787b3;
    ram[617] = 32'h40f707b3;
    ram[618] = 32'hd80306e3;
    ram[619] = 32'h267d7b3;
    ram[620] = 32'h1737;
    ram[621] = 32'hff470713;
    ram[622] = 32'hd6f77ee3;
    ram[623] = 32'h10737;
    ram[624] = 32'hff470713;
    ram[625] = 32'h4f76663;
    ram[626] = 32'h42423;
    ram[627] = 32'h2042823;
    ram[628] = 32'h513;
    ram[629] = 32'hd61ff06f;
    ram[630] = 32'h42e23;
    ram[631] = 32'he1dff06f;
    ram[632] = 32'h6b44783;
    ram[633] = 32'h6a44803;
    ram[634] = 32'h1879793;
    ram[635] = 32'h1081813;
    ram[636] = 32'h10787b3;
    ram[637] = 32'h6844803;
    ram[638] = 32'h10787b3;
    ram[639] = 32'h6944803;
    ram[640] = 32'h881813;
    ram[641] = 32'h10787b3;
    ram[642] = 32'h2f42023;
    ram[643] = 32'he79ff06f;
    ram[644] = 32'h100793;
    ram[645] = 32'h2f42823;
    ram[646] = 32'hfb9ff06f;
    ram[647] = 32'h54783;
    ram[648] = 32'hffe58593;
    ram[649] = 32'h2f585b3;
    ram[650] = 32'h452783;
    ram[651] = 32'hf585b3;
    ram[652] = 32'h3052783;
    ram[653] = 32'h79863;
    ram[654] = 32'h2855783;
    ram[655] = 32'h4047d793;
    ram[656] = 32'hf585b3;
    ram[657] = 32'h58513;
    ram[658] = 32'h8067;
    ram[659] = 32'h3452303;
    ram[660] = 32'h58793;
    ram[661] = 32'h78513;
    ram[662] = 32'h60593;
    ram[663] = 32'h68613;
    ram[664] = 32'h30067;
    ram[665] = 32'h3052783;
    ram[666] = 32'hfe010113;
    ram[667] = 32'h812c23;
    ram[668] = 32'h912a23;
    ram[669] = 32'h1312623;
    ram[670] = 32'h112e23;
    ram[671] = 32'h1212823;
    ram[672] = 32'h1412423;
    ram[673] = 32'h1512223;
    ram[674] = 32'h50493;
    ram[675] = 32'h60413;
    ram[676] = 32'h68993;
    ram[677] = 32'h6079e63;
    ram[678] = 32'h6059c63;
    ram[679] = 32'h1052783;
    ram[680] = 32'h2f66663;
    ram[681] = 32'h513;
    ram[682] = 32'h1c12083;
    ram[683] = 32'h1812403;
    ram[684] = 32'h1412483;
    ram[685] = 32'h1012903;
    ram[686] = 32'hc12983;
    ram[687] = 32'h812a03;
    ram[688] = 32'h412a83;
    ram[689] = 32'h2010113;
    ram[690] = 32'h8067;
    ram[691] = 32'h1c52503;
    ram[692] = 32'hc4a603;
    ram[693] = 32'hc50533;
    ram[694] = 32'ha40533;
    ram[695] = 32'h6098863;
    ram[696] = 32'h344a303;
    ram[697] = 32'h100613;
    ram[698] = 32'h98593;
    ram[699] = 32'h1812403;
    ram[700] = 32'h1c12083;
    ram[701] = 32'h1412483;
    ram[702] = 32'h1012903;
    ram[703] = 32'hc12983;
    ram[704] = 32'h812a03;
    ram[705] = 32'h412a83;
    ram[706] = 32'h2010113;
    ram[707] = 32'h30067;
    ram[708] = 32'h4ca03;
    ram[709] = 32'h913;
    ram[710] = 32'h3445ab3;
    ram[711] = 32'h1591e63;
    ram[712] = 32'hfff00793;
    ram[713] = 32'hf8f580e3;
    ram[714] = 32'h48513;
    ram[715] = 32'hef1ff0ef;
    ram[716] = 32'h3447433;
    ram[717] = 32'hfa5ff06f;
    ram[718] = 32'h48513;
    ram[719] = 32'hb8010ef;
    ram[720] = 32'h50593;
    ram[721] = 32'h190913;
    ram[722] = 32'hfd5ff06f;
    ram[723] = 32'h2444a783;
    ram[724] = 32'ha78c63;
    ram[725] = 32'h24a4a223;
    ram[726] = 32'h344a303;
    ram[727] = 32'h100613;
    ram[728] = 32'h4448593;
    ram[729] = 32'hf89ff06f;
    ram[730] = 32'h100513;
    ram[731] = 32'hf3dff06f;
    ram[732] = 32'h852503;
    ram[733] = 32'h8067;
    ram[734] = 32'hfb010113;
    ram[735] = 32'h5212023;
    ram[736] = 32'h3512a23;
    ram[737] = 32'h50913;
    ram[738] = 32'h58a93;
    ram[739] = 32'hc10513;
    ram[740] = 32'h100593;
    ram[741] = 32'h4912223;
    ram[742] = 32'h3312e23;
    ram[743] = 32'h3612823;
    ram[744] = 32'h3712623;
    ram[745] = 32'h3812423;
    ram[746] = 32'h3912223;
    ram[747] = 32'h4112623;
    ram[748] = 32'h4812423;
    ram[749] = 32'h3412c23;
    ram[750] = 32'h60b13;
    ram[751] = 32'h68b93;
    ram[752] = 32'h493;
    ram[753] = 32'h5dd000ef;
    ram[754] = 32'h24490c13;
    ram[755] = 32'h2000993;
    ram[756] = 32'h2000c93;
    ram[757] = 32'h693;
    ram[758] = 32'h48613;
    ram[759] = 32'ha8593;
    ram[760] = 32'h90513;
    ram[761] = 32'he81ff0ef;
    ram[762] = 32'h10050063;
    ram[763] = 32'h4490413;
    ram[764] = 32'h2e00a13;
    ram[765] = 32'h40513;
    ram[766] = 32'h5b1000ef;
    ram[767] = 32'hc050e63;
    ram[768] = 32'h12823;
    ram[769] = 32'h12a23;
    ram[770] = 32'h12c23;
    ram[771] = 32'h10e23;
    ram[772] = 32'h1010713;
    ram[773] = 32'h840693;
    ram[774] = 32'h40793;
    ram[775] = 32'h7c603;
    ram[776] = 32'h178793;
    ram[777] = 32'h170713;
    ram[778] = 32'hfec70fa3;
    ram[779] = 32'hfef698e3;
    ram[780] = 32'h844783;
    ram[781] = 32'h944683;
    ram[782] = 32'h100713;
    ram[783] = 32'hf10ca3;
    ram[784] = 32'hd10d23;
    ram[785] = 32'h1369663;
    ram[786] = 32'hfe078793;
    ram[787] = 32'hf03733;
    ram[788] = 32'ha44783;
    ram[789] = 32'hf10da3;
    ram[790] = 32'h1379463;
    ram[791] = 32'h6070463;
    ram[792] = 32'h1014783;
    ram[793] = 32'h7478063;
    ram[794] = 32'h1410c23;
    ram[795] = 32'hb0593;
    ram[796] = 32'h1010513;
    ram[797] = 32'h348000ef;
    ram[798] = 32'h4050a63;
    ram[799] = 32'h2000613;
    ram[800] = 32'h40593;
    ram[801] = 32'hb8513;
    ram[802] = 32'h98010ef;
    ram[803] = 32'h100513;
    ram[804] = 32'h4c12083;
    ram[805] = 32'h4812403;
    ram[806] = 32'h4412483;
    ram[807] = 32'h4012903;
    ram[808] = 32'h3c12983;
    ram[809] = 32'h3812a03;
    ram[810] = 32'h3412a83;
    ram[811] = 32'h3012b03;
    ram[812] = 32'h2c12b83;
    ram[813] = 32'h2812c03;
    ram[814] = 32'h2412c83;
    ram[815] = 32'h5010113;
    ram[816] = 32'h8067;
    ram[817] = 32'h1910c23;
    ram[818] = 32'hfa5ff06f;
    ram[819] = 32'h593;
    ram[820] = 32'hc10513;
    ram[821] = 32'h4cd000ef;
    ram[822] = 32'h2040413;
    ram[823] = 32'hf08c1ce3;
    ram[824] = 32'h148493;
    ram[825] = 32'hef1ff06f;
    ram[826] = 32'h513;
    ram[827] = 32'hfa5ff06f;
    ram[828] = 32'hc50633;
    ram[829] = 32'h1900313;
    ram[830] = 32'hc51863;
    ram[831] = 32'h793;
    ram[832] = 32'h78513;
    ram[833] = 32'h8067;
    ram[834] = 32'h54683;
    ram[835] = 32'h5c703;
    ram[836] = 32'hfbf68813;
    ram[837] = 32'hff87813;
    ram[838] = 32'h68793;
    ram[839] = 32'h1036663;
    ram[840] = 32'h2068793;
    ram[841] = 32'hff7f793;
    ram[842] = 32'hfbf70893;
    ram[843] = 32'hff8f893;
    ram[844] = 32'h70813;
    ram[845] = 32'h1136663;
    ram[846] = 32'h2070813;
    ram[847] = 32'hff87813;
    ram[848] = 32'h410787b3;
    ram[849] = 32'hfa079ee3;
    ram[850] = 32'hfa068ce3;
    ram[851] = 32'hfa070ae3;
    ram[852] = 32'h150513;
    ram[853] = 32'h158593;
    ram[854] = 32'hfa1ff06f;
    ram[855] = 32'h50793;
    ram[856] = 32'hfff00713;
    ram[857] = 32'h2e00613;
    ram[858] = 32'h7c683;
    ram[859] = 32'h69663;
    ram[860] = 32'h70513;
    ram[861] = 32'h8067;
    ram[862] = 32'hc69463;
    ram[863] = 32'h40a78733;
    ram[864] = 32'h178793;
    ram[865] = 32'hfe5ff06f;
    ram[866] = 32'h50793;
    ram[867] = 32'h6050463;
    ram[868] = 32'h54703;
    ram[869] = 32'h2f00693;
    ram[870] = 32'hd71863;
    ram[871] = 32'h150793;
    ram[872] = 32'h513;
    ram[873] = 32'h400006f;
    ram[874] = 32'h154683;
    ram[875] = 32'h3a00713;
    ram[876] = 32'he68a63;
    ram[877] = 32'h254683;
    ram[878] = 32'h5c00713;
    ram[879] = 32'hfff00513;
    ram[880] = 32'h2e69c63;
    ram[881] = 32'h378793;
    ram[882] = 32'h5c00713;
    ram[883] = 32'hfd5ff06f;
    ram[884] = 32'h178793;
    ram[885] = 32'he68663;
    ram[886] = 32'h7c683;
    ram[887] = 32'hfe069ae3;
    ram[888] = 32'h150513;
    ram[889] = 32'h7c683;
    ram[890] = 32'hfe0698e3;
    ram[891] = 32'hfff50513;
    ram[892] = 32'h8067;
    ram[893] = 32'hfff00513;
    ram[894] = 32'h8067;
    ram[895] = 32'hfff00793;
    ram[896] = 32'he050263;
    ram[897] = 32'hed05063;
    ram[898] = 32'hfe010113;
    ram[899] = 32'h812c23;
    ram[900] = 32'h112e23;
    ram[901] = 32'h912a23;
    ram[902] = 32'h1212823;
    ram[903] = 32'h1312623;
    ram[904] = 32'h1412423;
    ram[905] = 32'h54983;
    ram[906] = 32'h2f00793;
    ram[907] = 32'h150413;
    ram[908] = 32'h2f98463;
    ram[909] = 32'h154703;
    ram[910] = 32'h3a00793;
    ram[911] = 32'hf70a63;
    ram[912] = 32'h254803;
    ram[913] = 32'h5c00713;
    ram[914] = 32'hfff00793;
    ram[915] = 32'h4e81663;
    ram[916] = 32'h350413;
    ram[917] = 32'h5c00993;
    ram[918] = 32'h40513;
    ram[919] = 32'h68493;
    ram[920] = 32'h60913;
    ram[921] = 32'h58a13;
    ram[922] = 32'h69d000ef;
    ram[923] = 32'h40793;
    ram[924] = 32'h713;
    ram[925] = 32'h613;
    ram[926] = 32'hfff48693;
    ram[927] = 32'h408785b3;
    ram[928] = 32'he90833;
    ram[929] = 32'h2a5cc63;
    ram[930] = 32'h80023;
    ram[931] = 32'h94783;
    ram[932] = 32'h17b793;
    ram[933] = 32'h40f007b3;
    ram[934] = 32'h1c12083;
    ram[935] = 32'h1812403;
    ram[936] = 32'h1412483;
    ram[937] = 32'h1012903;
    ram[938] = 32'hc12983;
    ram[939] = 32'h812a03;
    ram[940] = 32'h78513;
    ram[941] = 32'h2010113;
    ram[942] = 32'h8067;
    ram[943] = 32'h7c583;
    ram[944] = 32'h1359863;
    ram[945] = 32'h160613;
    ram[946] = 32'h178793;
    ram[947] = 32'hfb1ff06f;
    ram[948] = 32'hff461ce3;
    ram[949] = 32'hfed75ae3;
    ram[950] = 32'h170713;
    ram[951] = 32'hb80023;
    ram[952] = 32'hfe9ff06f;
    ram[953] = 32'h78513;
    ram[954] = 32'h8067;
    ram[955] = 32'hfd010113;
    ram[956] = 32'h2912223;
    ram[957] = 32'h3212023;
    ram[958] = 32'h1312e23;
    ram[959] = 32'h1412c23;
    ram[960] = 32'he12623;
    ram[961] = 32'h2112623;
    ram[962] = 32'h2812423;
    ram[963] = 32'h50913;
    ram[964] = 32'h58493;
    ram[965] = 32'h60993;
    ram[966] = 32'h68a13;
    ram[967] = 32'he6dff0ef;
    ram[968] = 32'hfff00793;
    ram[969] = 32'hc12703;
    ram[970] = 32'h2f51663;
    ram[971] = 32'hfff00413;
    ram[972] = 32'h40513;
    ram[973] = 32'h2c12083;
    ram[974] = 32'h2812403;
    ram[975] = 32'h2412483;
    ram[976] = 32'h2012903;
    ram[977] = 32'h1c12983;
    ram[978] = 32'h1812a03;
    ram[979] = 32'h3010113;
    ram[980] = 32'h8067;
    ram[981] = 32'h50413;
    ram[982] = 32'h50593;
    ram[983] = 32'h70693;
    ram[984] = 32'ha0613;
    ram[985] = 32'h90513;
    ram[986] = 32'he95ff0ef;
    ram[987] = 32'hfc0510e3;
    ram[988] = 32'h41663;
    ram[989] = 32'h48023;
    ram[990] = 32'hfb9ff06f;
    ram[991] = 32'h90513;
    ram[992] = 32'h585000ef;
    ram[993] = 32'h50413;
    ram[994] = 32'ha0513;
    ram[995] = 32'h579000ef;
    ram[996] = 32'h40a40433;
    ram[997] = 32'h89d463;
    ram[998] = 32'h98413;
    ram[999] = 32'h40613;
    ram[1000] = 32'h90593;
    ram[1001] = 32'h848433;
    ram[1002] = 32'h48513;
    ram[1003] = 32'h575000ef;
    ram[1004] = 32'hfe040fa3;
    ram[1005] = 32'h413;
    ram[1006] = 32'hf79ff06f;
    ram[1007] = 32'hfd010113;
    ram[1008] = 32'h2112623;
    ram[1009] = 32'h2812423;
    ram[1010] = 32'h2912223;
    ram[1011] = 32'h3212023;
    ram[1012] = 32'h1312e23;
    ram[1013] = 32'h58913;
    ram[1014] = 32'h1412c23;
    ram[1015] = 32'h1512a23;
    ram[1016] = 32'h1612823;
    ram[1017] = 32'h50a13;
    ram[1018] = 32'hd75ff0ef;
    ram[1019] = 32'h50493;
    ram[1020] = 32'h90513;
    ram[1021] = 32'hd69ff0ef;
    ram[1022] = 32'hfff00793;
    ram[1023] = 32'h50413;
    ram[1024] = 32'h993;
    ram[1025] = 32'h8f49c63;
    ram[1026] = 32'hc951c63;
    ram[1027] = 32'ha0513;
    ram[1028] = 32'h4f5000ef;
    ram[1029] = 32'h50493;
    ram[1030] = 32'h90513;
    ram[1031] = 32'h4e9000ef;
    ram[1032] = 32'h50413;
    ram[1033] = 32'hfff48793;
    ram[1034] = 32'hfa07b3;
    ram[1035] = 32'h40f486b3;
    ram[1036] = 32'h2000613;
    ram[1037] = 32'hd78733;
    ram[1038] = 32'h70663;
    ram[1039] = 32'h7c703;
    ram[1040] = 32'h4c70263;
    ram[1041] = 32'hfff40793;
    ram[1042] = 32'hf907b3;
    ram[1043] = 32'h40f406b3;
    ram[1044] = 32'h2000613;
    ram[1045] = 32'hd78733;
    ram[1046] = 32'h70663;
    ram[1047] = 32'h7c703;
    ram[1048] = 32'h2c70863;
    ram[1049] = 32'h993;
    ram[1050] = 32'h6941c63;
    ram[1051] = 32'h40613;
    ram[1052] = 32'h90593;
    ram[1053] = 32'ha0513;
    ram[1054] = 32'hc79ff0ef;
    ram[1055] = 32'h153993;
    ram[1056] = 32'h600006f;
    ram[1057] = 32'h414784b3;
    ram[1058] = 32'hfff78793;
    ram[1059] = 32'hfa9ff06f;
    ram[1060] = 32'h41278433;
    ram[1061] = 32'hfff78793;
    ram[1062] = 32'hfbdff06f;
    ram[1063] = 32'h4f50263;
    ram[1064] = 32'h148a93;
    ram[1065] = 32'h15a0ab3;
    ram[1066] = 32'h140b13;
    ram[1067] = 32'ha8513;
    ram[1068] = 32'h455000ef;
    ram[1069] = 32'h1690b33;
    ram[1070] = 32'ha12623;
    ram[1071] = 32'hb0513;
    ram[1072] = 32'h445000ef;
    ram[1073] = 32'hc12603;
    ram[1074] = 32'h993;
    ram[1075] = 32'ha61a63;
    ram[1076] = 32'hb0593;
    ram[1077] = 32'ha8513;
    ram[1078] = 32'hc19ff0ef;
    ram[1079] = 32'hf40504e3;
    ram[1080] = 32'h2c12083;
    ram[1081] = 32'h2812403;
    ram[1082] = 32'h98513;
    ram[1083] = 32'h2412483;
    ram[1084] = 32'h2012903;
    ram[1085] = 32'h1c12983;
    ram[1086] = 32'h1812a03;
    ram[1087] = 32'h1412a83;
    ram[1088] = 32'h1012b03;
    ram[1089] = 32'h3010113;
    ram[1090] = 32'h8067;
    ram[1091] = 32'hfc010113;
    ram[1092] = 32'h2812c23;
    ram[1093] = 32'h82000437;
    ram[1094] = 32'h46444783;
    ram[1095] = 32'h3512223;
    ram[1096] = 32'h3212823;
    ram[1097] = 32'h2f5fab3;
    ram[1098] = 32'h3412423;
    ram[1099] = 32'h3612023;
    ram[1100] = 32'h1712e23;
    ram[1101] = 32'h2112e23;
    ram[1102] = 32'h2912a23;
    ram[1103] = 32'h3312623;
    ram[1104] = 32'h50913;
    ram[1105] = 32'h60b93;
    ram[1106] = 32'h1568733;
    ram[1107] = 32'h2f5da33;
    ram[1108] = 32'h41578b33;
    ram[1109] = 32'he7e463;
    ram[1110] = 32'h68b13;
    ram[1111] = 32'h22892983;
    ram[1112] = 32'h7499463;
    ram[1113] = 32'h22c92483;
    ram[1114] = 32'hfff00793;
    ram[1115] = 32'h2f48463;
    ram[1116] = 32'h48593;
    ram[1117] = 32'h46440513;
    ram[1118] = 32'h8a5ff0ef;
    ram[1119] = 32'h15505b3;
    ram[1120] = 32'hb0693;
    ram[1121] = 32'hb8613;
    ram[1122] = 32'h46440513;
    ram[1123] = 32'h8c1ff0ef;
    ram[1124] = 32'h51463;
    ram[1125] = 32'hb13;
    ram[1126] = 32'h3c12083;
    ram[1127] = 32'h3812403;
    ram[1128] = 32'hb0513;
    ram[1129] = 32'h3412483;
    ram[1130] = 32'h3012903;
    ram[1131] = 32'h2c12983;
    ram[1132] = 32'h2812a03;
    ram[1133] = 32'h2412a83;
    ram[1134] = 32'h2012b03;
    ram[1135] = 32'h1c12b83;
    ram[1136] = 32'h4010113;
    ram[1137] = 32'h8067;
    ram[1138] = 32'h20a0463;
    ram[1139] = 32'h198793;
    ram[1140] = 32'h3479063;
    ram[1141] = 32'h22c92483;
    ram[1142] = 32'h349e263;
    ram[1143] = 32'hfff00793;
    ram[1144] = 32'hfaf48ae3;
    ram[1145] = 32'h22992623;
    ram[1146] = 32'h23492423;
    ram[1147] = 32'hf85ff06f;
    ram[1148] = 32'h492483;
    ram[1149] = 32'h993;
    ram[1150] = 32'hfe1ff06f;
    ram[1151] = 32'hc10693;
    ram[1152] = 32'h98613;
    ram[1153] = 32'h90593;
    ram[1154] = 32'h46440513;
    ram[1155] = 32'hce4ff0ef;
    ram[1156] = 32'h2051463;
    ram[1157] = 32'h48593;
    ram[1158] = 32'h46440513;
    ram[1159] = 32'h1d9000ef;
    ram[1160] = 32'h50693;
    ram[1161] = 32'ha12623;
    ram[1162] = 32'h98613;
    ram[1163] = 32'h90593;
    ram[1164] = 32'h46440513;
    ram[1165] = 32'hcc4ff0ef;
    ram[1166] = 32'hc12483;
    ram[1167] = 32'h198993;
    ram[1168] = 32'hf99ff06f;
    ram[1169] = 32'h452783;
    ram[1170] = 32'h4079463;
    ram[1171] = 32'h52783;
    ram[1172] = 32'h79c63;
    ram[1173] = 32'hb52023;
    ram[1174] = 32'hb52223;
    ram[1175] = 32'h5a023;
    ram[1176] = 32'h5a223;
    ram[1177] = 32'h8067;
    ram[1178] = 32'h7a703;
    ram[1179] = 32'hf5a223;
    ram[1180] = 32'he5a023;
    ram[1181] = 32'h7a703;
    ram[1182] = 32'h71863;
    ram[1183] = 32'hb52023;
    ram[1184] = 32'hb7a023;
    ram[1185] = 32'h8067;
    ram[1186] = 32'hb72223;
    ram[1187] = 32'hff5ff06f;
    ram[1188] = 32'h47a703;
    ram[1189] = 32'hf5a023;
    ram[1190] = 32'he5a223;
    ram[1191] = 32'h47a703;
    ram[1192] = 32'h71863;
    ram[1193] = 32'hb52223;
    ram[1194] = 32'hb7a223;
    ram[1195] = 32'h8067;
    ram[1196] = 32'hb72023;
    ram[1197] = 32'hff5ff06f;
    ram[1198] = 32'h43c52783;
    ram[1199] = 32'h43c50593;
    ram[1200] = 32'h44052703;
    ram[1201] = 32'h2079463;
    ram[1202] = 32'h820016b7;
    ram[1203] = 32'h8ee6a223;
    ram[1204] = 32'h44052703;
    ram[1205] = 32'h2071063;
    ram[1206] = 32'h82001737;
    ram[1207] = 32'h8ef72423;
    ram[1208] = 32'h82001537;
    ram[1209] = 32'h8dc50513;
    ram[1210] = 32'hf5dff06f;
    ram[1211] = 32'he7a223;
    ram[1212] = 32'hfe1ff06f;
    ram[1213] = 32'hf72023;
    ram[1214] = 32'hfe9ff06f;
    ram[1215] = 32'hea010113;
    ram[1216] = 32'h820017b7;
    ram[1217] = 32'h14912a23;
    ram[1218] = 32'h8dc7a483;
    ram[1219] = 32'h14112e23;
    ram[1220] = 32'h14812c23;
    ram[1221] = 32'h15212823;
    ram[1222] = 32'h15312623;
    ram[1223] = 32'h15412423;
    ram[1224] = 32'h15512223;
    ram[1225] = 32'h15612023;
    ram[1226] = 32'h13712e23;
    ram[1227] = 32'h13812c23;
    ram[1228] = 32'h49663;
    ram[1229] = 32'h413;
    ram[1230] = 32'h1ac0006f;
    ram[1231] = 32'h4a703;
    ram[1232] = 32'h8dc78793;
    ram[1233] = 32'h44a683;
    ram[1234] = 32'h8071663;
    ram[1235] = 32'hd7a023;
    ram[1236] = 32'h44a683;
    ram[1237] = 32'h8069463;
    ram[1238] = 32'he7a223;
    ram[1239] = 32'h50913;
    ram[1240] = 32'h82001537;
    ram[1241] = 32'h8e450993;
    ram[1242] = 32'h48593;
    ram[1243] = 32'h8e450513;
    ram[1244] = 32'hed5ff0ef;
    ram[1245] = 32'h43c00793;
    ram[1246] = 32'hbc448413;
    ram[1247] = 32'hfaf48ce3;
    ram[1248] = 32'hbd848a13;
    ram[1249] = 32'h10400613;
    ram[1250] = 32'h593;
    ram[1251] = 32'ha0513;
    ram[1252] = 32'h1b5000ef;
    ram[1253] = 32'hcdc48a93;
    ram[1254] = 32'h10400613;
    ram[1255] = 32'h593;
    ram[1256] = 32'ha8513;
    ram[1257] = 32'h1a1000ef;
    ram[1258] = 32'h10400713;
    ram[1259] = 32'ha8693;
    ram[1260] = 32'h10400613;
    ram[1261] = 32'ha0593;
    ram[1262] = 32'h90513;
    ram[1263] = 32'hb31ff0ef;
    ram[1264] = 32'hfff00793;
    ram[1265] = 32'h2f51063;
    ram[1266] = 32'h40513;
    ram[1267] = 32'heedff0ef;
    ram[1268] = 32'hf65ff06f;
    ram[1269] = 32'hd72223;
    ram[1270] = 32'hf79ff06f;
    ram[1271] = 32'he6a023;
    ram[1272] = 32'hf7dff06f;
    ram[1273] = 32'h9a903;
    ram[1274] = 32'h2091e63;
    ram[1275] = 32'h1444783;
    ram[1276] = 32'h820009b7;
    ram[1277] = 32'h6078263;
    ram[1278] = 32'h46498513;
    ram[1279] = 32'hf74ff0ef;
    ram[1280] = 32'h50913;
    ram[1281] = 32'ha0513;
    ram[1282] = 32'h981ff0ef;
    ram[1283] = 32'h50b93;
    ram[1284] = 32'hb13;
    ram[1285] = 32'hfff00c13;
    ram[1286] = 32'h116bd063;
    ram[1287] = 32'hbd24a223;
    ram[1288] = 32'h440006f;
    ram[1289] = 32'hbc490793;
    ram[1290] = 32'hf41663;
    ram[1291] = 32'h492903;
    ram[1292] = 32'hfb9ff06f;
    ram[1293] = 32'ha0593;
    ram[1294] = 32'hbd890513;
    ram[1295] = 32'hb81ff0ef;
    ram[1296] = 32'hfe0506e3;
    ram[1297] = 32'ha8593;
    ram[1298] = 32'hcdc90513;
    ram[1299] = 32'hb71ff0ef;
    ram[1300] = 32'hfc050ee3;
    ram[1301] = 32'hf75ff06f;
    ram[1302] = 32'h46498513;
    ram[1303] = 32'hf14ff0ef;
    ram[1304] = 32'hbca4a223;
    ram[1305] = 32'hbc44a583;
    ram[1306] = 32'h2c10693;
    ram[1307] = 32'ha8613;
    ram[1308] = 32'h46498513;
    ram[1309] = 32'hf04ff0ef;
    ram[1310] = 32'hf40508e3;
    ram[1311] = 32'h2c10513;
    ram[1312] = 32'h574000ef;
    ram[1313] = 32'hf40502e3;
    ram[1314] = 32'hb00613;
    ram[1315] = 32'h2c10593;
    ram[1316] = 32'h21c40513;
    ram[1317] = 32'h8d000ef;
    ram[1318] = 32'h4812783;
    ram[1319] = 32'h42423;
    ram[1320] = 32'h40593;
    ram[1321] = 32'hf42623;
    ram[1322] = 32'h4015783;
    ram[1323] = 32'h4615703;
    ram[1324] = 32'h46498513;
    ram[1325] = 32'h1079793;
    ram[1326] = 32'he787b3;
    ram[1327] = 32'hf42223;
    ram[1328] = 32'hfff00793;
    ram[1329] = 32'h42f42823;
    ram[1330] = 32'h42042a23;
    ram[1331] = 32'h42823;
    ram[1332] = 32'h22f42423;
    ram[1333] = 32'h22f42623;
    ram[1334] = 32'ha10ff0ef;
    ram[1335] = 32'h46498513;
    ram[1336] = 32'h6bc000ef;
    ram[1337] = 32'h40513;
    ram[1338] = 32'h15c12083;
    ram[1339] = 32'h15812403;
    ram[1340] = 32'h15412483;
    ram[1341] = 32'h15012903;
    ram[1342] = 32'h14c12983;
    ram[1343] = 32'h14812a03;
    ram[1344] = 32'h14412a83;
    ram[1345] = 32'h14012b03;
    ram[1346] = 32'h13c12b83;
    ram[1347] = 32'h13812c03;
    ram[1348] = 32'h16010113;
    ram[1349] = 32'h8067;
    ram[1350] = 32'h10400693;
    ram[1351] = 32'h2c10613;
    ram[1352] = 32'hb0593;
    ram[1353] = 32'ha0513;
    ram[1354] = 32'h8d5ff0ef;
    ram[1355] = 32'he9850ee3;
    ram[1356] = 32'hc10693;
    ram[1357] = 32'h2c10613;
    ram[1358] = 32'h90593;
    ram[1359] = 32'h46498513;
    ram[1360] = 32'he38ff0ef;
    ram[1361] = 32'he80502e3;
    ram[1362] = 32'hc10513;
    ram[1363] = 32'h498000ef;
    ram[1364] = 32'he6050ce3;
    ram[1365] = 32'h2015903;
    ram[1366] = 32'h2615783;
    ram[1367] = 32'h1b0b13;
    ram[1368] = 32'h1091913;
    ram[1369] = 32'hf90933;
    ram[1370] = 32'heb1ff06f;
    ram[1371] = 32'hff010113;
    ram[1372] = 32'h82001537;
    ram[1373] = 32'h112623;
    ram[1374] = 32'h8dc50793;
    ram[1375] = 32'h7a223;
    ram[1376] = 32'h7a023;
    ram[1377] = 32'h820005b7;
    ram[1378] = 32'h820017b7;
    ram[1379] = 32'h8e478793;
    ram[1380] = 32'h45c58593;
    ram[1381] = 32'h8dc50513;
    ram[1382] = 32'h7a223;
    ram[1383] = 32'h7a023;
    ram[1384] = 32'hca5ff0ef;
    ram[1385] = 32'hc12083;
    ram[1386] = 32'h820017b7;
    ram[1387] = 32'h100713;
    ram[1388] = 32'h8ce7aa23;
    ram[1389] = 32'h1010113;
    ram[1390] = 32'h8067;
    ram[1391] = 32'h820017b7;
    ram[1392] = 32'h8d47a783;
    ram[1393] = 32'hfe010113;
    ram[1394] = 32'h112e23;
    ram[1395] = 32'h79c63;
    ram[1396] = 32'hb12623;
    ram[1397] = 32'ha12423;
    ram[1398] = 32'hf95ff0ef;
    ram[1399] = 32'hc12583;
    ram[1400] = 32'h812503;
    ram[1401] = 32'h820007b7;
    ram[1402] = 32'h46478713;
    ram[1403] = 32'h2a72a23;
    ram[1404] = 32'h46478513;
    ram[1405] = 32'h2b72c23;
    ram[1406] = 32'h908ff0ef;
    ram[1407] = 32'h51863;
    ram[1408] = 32'h820017b7;
    ram[1409] = 32'h100713;
    ram[1410] = 32'h8ce7ac23;
    ram[1411] = 32'h1c12083;
    ram[1412] = 32'h2010113;
    ram[1413] = 32'h8067;
    ram[1414] = 32'h820017b7;
    ram[1415] = 32'h8d47a783;
    ram[1416] = 32'hfe010113;
    ram[1417] = 32'h912a23;
    ram[1418] = 32'h1212823;
    ram[1419] = 32'h112e23;
    ram[1420] = 32'h812c23;
    ram[1421] = 32'h50913;
    ram[1422] = 32'h58493;
    ram[1423] = 32'h79463;
    ram[1424] = 32'hf2dff0ef;
    ram[1425] = 32'h820017b7;
    ram[1426] = 32'h8d87a783;
    ram[1427] = 32'h513;
    ram[1428] = 32'h8078a63;
    ram[1429] = 32'h8090863;
    ram[1430] = 32'h8048663;
    ram[1431] = 32'h48513;
    ram[1432] = 32'h6a4000ef;
    ram[1433] = 32'h48713;
    ram[1434] = 32'h413;
    ram[1435] = 32'h5700693;
    ram[1436] = 32'h6200613;
    ram[1437] = 32'h7200813;
    ram[1438] = 32'h7700893;
    ram[1439] = 32'h6100313;
    ram[1440] = 32'h4100593;
    ram[1441] = 32'h4200e13;
    ram[1442] = 32'h5200e93;
    ram[1443] = 32'h2b00f13;
    ram[1444] = 32'h409707b3;
    ram[1445] = 32'h6a7c463;
    ram[1446] = 32'h820007b7;
    ram[1447] = 32'h46478713;
    ram[1448] = 32'h3c72703;
    ram[1449] = 32'h46478493;
    ram[1450] = 32'h70463;
    ram[1451] = 32'h700e7;
    ram[1452] = 32'h147793;
    ram[1453] = 32'h513;
    ram[1454] = 32'h78c63;
    ram[1455] = 32'h90513;
    ram[1456] = 32'hc3dff0ef;
    ram[1457] = 32'h50663;
    ram[1458] = 32'hfd947413;
    ram[1459] = 32'h42850c23;
    ram[1460] = 32'h404a783;
    ram[1461] = 32'h78863;
    ram[1462] = 32'ha12623;
    ram[1463] = 32'h780e7;
    ram[1464] = 32'hc12503;
    ram[1465] = 32'h1c12083;
    ram[1466] = 32'h1812403;
    ram[1467] = 32'h1412483;
    ram[1468] = 32'h1012903;
    ram[1469] = 32'h2010113;
    ram[1470] = 32'h8067;
    ram[1471] = 32'h74783;
    ram[1472] = 32'h4d78463;
    ram[1473] = 32'h2f6e463;
    ram[1474] = 32'h2b78863;
    ram[1475] = 32'hf5e863;
    ram[1476] = 32'h5e78063;
    ram[1477] = 32'h170713;
    ram[1478] = 32'hf79ff06f;
    ram[1479] = 32'h7c78263;
    ram[1480] = 32'hffd79ae3;
    ram[1481] = 32'h146413;
    ram[1482] = 32'hfedff06f;
    ram[1483] = 32'h4c78a63;
    ram[1484] = 32'hf66863;
    ram[1485] = 32'hfe6790e3;
    ram[1486] = 32'h2646413;
    ram[1487] = 32'hfd9ff06f;
    ram[1488] = 32'hff0782e3;
    ram[1489] = 32'hfd1798e3;
    ram[1490] = 32'h3246413;
    ram[1491] = 32'hfc9ff06f;
    ram[1492] = 32'h147793;
    ram[1493] = 32'h78663;
    ram[1494] = 32'h246413;
    ram[1495] = 32'hfb9ff06f;
    ram[1496] = 32'h247793;
    ram[1497] = 32'h78663;
    ram[1498] = 32'h3146413;
    ram[1499] = 32'hfa9ff06f;
    ram[1500] = 32'h447793;
    ram[1501] = 32'hfa0780e3;
    ram[1502] = 32'h2746413;
    ram[1503] = 32'hf99ff06f;
    ram[1504] = 32'h846413;
    ram[1505] = 32'hf91ff06f;
    ram[1506] = 32'h820017b7;
    ram[1507] = 32'h8d47a783;
    ram[1508] = 32'hff010113;
    ram[1509] = 32'h812423;
    ram[1510] = 32'h112623;
    ram[1511] = 32'h912223;
    ram[1512] = 32'h1212023;
    ram[1513] = 32'h50413;
    ram[1514] = 32'h79463;
    ram[1515] = 32'hdc1ff0ef;
    ram[1516] = 32'h6040463;
    ram[1517] = 32'h820004b7;
    ram[1518] = 32'h46448793;
    ram[1519] = 32'h3c7a783;
    ram[1520] = 32'h46448913;
    ram[1521] = 32'h78463;
    ram[1522] = 32'h780e7;
    ram[1523] = 32'hfff00793;
    ram[1524] = 32'h42f42823;
    ram[1525] = 32'h40513;
    ram[1526] = 32'h42423;
    ram[1527] = 32'h42623;
    ram[1528] = 32'h42223;
    ram[1529] = 32'h42042a23;
    ram[1530] = 32'h42823;
    ram[1531] = 32'hacdff0ef;
    ram[1532] = 32'h46448513;
    ram[1533] = 32'h3a8000ef;
    ram[1534] = 32'h4092303;
    ram[1535] = 32'h30e63;
    ram[1536] = 32'h812403;
    ram[1537] = 32'hc12083;
    ram[1538] = 32'h412483;
    ram[1539] = 32'h12903;
    ram[1540] = 32'h1010113;
    ram[1541] = 32'h30067;
    ram[1542] = 32'hc12083;
    ram[1543] = 32'h812403;
    ram[1544] = 32'h412483;
    ram[1545] = 32'h12903;
    ram[1546] = 32'h1010113;
    ram[1547] = 32'h8067;
    ram[1548] = 32'h820017b7;
    ram[1549] = 32'h8d47a783;
    ram[1550] = 32'hfd010113;
    ram[1551] = 32'h2812423;
    ram[1552] = 32'h2912223;
    ram[1553] = 32'h1612823;
    ram[1554] = 32'h2112623;
    ram[1555] = 32'h3212023;
    ram[1556] = 32'h1312e23;
    ram[1557] = 32'h1412c23;
    ram[1558] = 32'h1512a23;
    ram[1559] = 32'h1712623;
    ram[1560] = 32'h1812423;
    ram[1561] = 32'h1912223;
    ram[1562] = 32'h50b13;
    ram[1563] = 32'h68493;
    ram[1564] = 32'h2c58433;
    ram[1565] = 32'h79463;
    ram[1566] = 32'hcf5ff0ef;
    ram[1567] = 32'h100b0e63;
    ram[1568] = 32'h10048c63;
    ram[1569] = 32'h4384c783;
    ram[1570] = 32'h17f793;
    ram[1571] = 32'h10078663;
    ram[1572] = 32'h2040e63;
    ram[1573] = 32'h84a583;
    ram[1574] = 32'hc4a783;
    ram[1575] = 32'hef5fe63;
    ram[1576] = 32'hb40733;
    ram[1577] = 32'h40a93;
    ram[1578] = 32'he7f463;
    ram[1579] = 32'h40b78ab3;
    ram[1580] = 32'h95d993;
    ram[1581] = 32'h1ff5f913;
    ram[1582] = 32'h413;
    ram[1583] = 32'h23048b93;
    ram[1584] = 32'h20000c13;
    ram[1585] = 32'h1ff00c93;
    ram[1586] = 32'h3544e63;
    ram[1587] = 32'h40513;
    ram[1588] = 32'h2c12083;
    ram[1589] = 32'h2812403;
    ram[1590] = 32'h2412483;
    ram[1591] = 32'h2012903;
    ram[1592] = 32'h1c12983;
    ram[1593] = 32'h1812a03;
    ram[1594] = 32'h1412a83;
    ram[1595] = 32'h1012b03;
    ram[1596] = 32'hc12b83;
    ram[1597] = 32'h812c03;
    ram[1598] = 32'h412c83;
    ram[1599] = 32'h3010113;
    ram[1600] = 32'h8067;
    ram[1601] = 32'h4091263;
    ram[1602] = 32'h408a86b3;
    ram[1603] = 32'h2dcde63;
    ram[1604] = 32'h4096d693;
    ram[1605] = 32'h8b0633;
    ram[1606] = 32'h98593;
    ram[1607] = 32'h48513;
    ram[1608] = 32'hfecff0ef;
    ram[1609] = 32'hfa0504e3;
    ram[1610] = 32'h951a13;
    ram[1611] = 32'ha989b3;
    ram[1612] = 32'h84a783;
    ram[1613] = 32'h1440433;
    ram[1614] = 32'h913;
    ram[1615] = 32'h1478a33;
    ram[1616] = 32'h144a423;
    ram[1617] = 32'hf85ff06f;
    ram[1618] = 32'h4304a783;
    ram[1619] = 32'h3378263;
    ram[1620] = 32'h100693;
    ram[1621] = 32'hb8613;
    ram[1622] = 32'h98593;
    ram[1623] = 32'h48513;
    ram[1624] = 32'hfacff0ef;
    ram[1625] = 32'hf60504e3;
    ram[1626] = 32'h4334a823;
    ram[1627] = 32'h4204aa23;
    ram[1628] = 32'h412c07b3;
    ram[1629] = 32'h408a8a33;
    ram[1630] = 32'h147d463;
    ram[1631] = 32'h78a13;
    ram[1632] = 32'ha0613;
    ram[1633] = 32'h12b85b3;
    ram[1634] = 32'h8b0533;
    ram[1635] = 32'h394000ef;
    ram[1636] = 32'h198993;
    ram[1637] = 32'hf9dff06f;
    ram[1638] = 32'hfff00413;
    ram[1639] = 32'hf31ff06f;
    ram[1640] = 32'h50023;
    ram[1641] = 32'h8067;
    ram[1642] = 32'hb54783;
    ram[1643] = 32'hf00713;
    ram[1644] = 32'h2e78663;
    ram[1645] = 32'h54703;
    ram[1646] = 32'h513;
    ram[1647] = 32'h2070263;
    ram[1648] = 32'he500693;
    ram[1649] = 32'hd70e63;
    ram[1650] = 32'h800713;
    ram[1651] = 32'he78a63;
    ram[1652] = 32'h67f793;
    ram[1653] = 32'h17b513;
    ram[1654] = 32'h8067;
    ram[1655] = 32'h513;
    ram[1656] = 32'h8067;
    ram[1657] = 32'hb54503;
    ram[1658] = 32'h455513;
    ram[1659] = 32'h157513;
    ram[1660] = 32'h8067;
    ram[1661] = 32'hb54503;
    ram[1662] = 32'h555513;
    ram[1663] = 32'h157513;
    ram[1664] = 32'h8067;
    ram[1665] = 32'h3852683;
    ram[1666] = 32'hff010113;
    ram[1667] = 32'h812423;
    ram[1668] = 32'h112623;
    ram[1669] = 32'h58413;
    ram[1670] = 32'h69e63;
    ram[1671] = 32'h20042223;
    ram[1672] = 32'h100513;
    ram[1673] = 32'hc12083;
    ram[1674] = 32'h812403;
    ram[1675] = 32'h1010113;
    ram[1676] = 32'h8067;
    ram[1677] = 32'h50713;
    ram[1678] = 32'h1472783;
    ram[1679] = 32'h2005a503;
    ram[1680] = 32'h2072703;
    ram[1681] = 32'h100613;
    ram[1682] = 32'h40f507b3;
    ram[1683] = 32'h178593;
    ram[1684] = 32'hb77463;
    ram[1685] = 32'h40f70633;
    ram[1686] = 32'h40593;
    ram[1687] = 32'h680e7;
    ram[1688] = 32'hfa051ee3;
    ram[1689] = 32'hfc1ff06f;
    ram[1690] = 32'hfe010113;
    ram[1691] = 32'h1212823;
    ram[1692] = 32'h25452903;
    ram[1693] = 32'h812c23;
    ram[1694] = 32'h112e23;
    ram[1695] = 32'h912a23;
    ram[1696] = 32'h1312623;
    ram[1697] = 32'h413;
    ram[1698] = 32'h6091a63;
    ram[1699] = 32'h25452783;
    ram[1700] = 32'h58493;
    ram[1701] = 32'h50993;
    ram[1702] = 32'h20f42623;
    ram[1703] = 32'h20442783;
    ram[1704] = 32'h24852a23;
    ram[1705] = 32'h78a63;
    ram[1706] = 32'h40593;
    ram[1707] = 32'h98513;
    ram[1708] = 32'hf55ff0ef;
    ram[1709] = 32'h2050463;
    ram[1710] = 32'h349a783;
    ram[1711] = 32'h20942023;
    ram[1712] = 32'h100613;
    ram[1713] = 32'h40593;
    ram[1714] = 32'h48513;
    ram[1715] = 32'h780e7;
    ram[1716] = 32'h6051063;
    ram[1717] = 32'hfff00793;
    ram[1718] = 32'h20f42023;
    ram[1719] = 32'h1c12083;
    ram[1720] = 32'h1812403;
    ram[1721] = 32'h90513;
    ram[1722] = 32'h1412483;
    ram[1723] = 32'h1012903;
    ram[1724] = 32'hc12983;
    ram[1725] = 32'h2010113;
    ram[1726] = 32'h8067;
    ram[1727] = 32'h20092783;
    ram[1728] = 32'hf5e663;
    ram[1729] = 32'h178713;
    ram[1730] = 32'h2e5ea63;
    ram[1731] = 32'h20c92783;
    ram[1732] = 32'h79663;
    ram[1733] = 32'h40a63;
    ram[1734] = 32'h20042623;
    ram[1735] = 32'h90413;
    ram[1736] = 32'h20c92903;
    ram[1737] = 32'hf65ff06f;
    ram[1738] = 32'h24052a23;
    ram[1739] = 32'hff1ff06f;
    ram[1740] = 32'h20842423;
    ram[1741] = 32'h40913;
    ram[1742] = 32'hfa5ff06f;
    ram[1743] = 32'h40f585b3;
    ram[1744] = 32'h959593;
    ram[1745] = 32'hb905b3;
    ram[1746] = 32'h20b92423;
    ram[1747] = 32'hf91ff06f;
    ram[1748] = 32'hff010113;
    ram[1749] = 32'h812423;
    ram[1750] = 32'h112623;
    ram[1751] = 32'hfff00793;
    ram[1752] = 32'h44f52c23;
    ram[1753] = 32'h25850793;
    ram[1754] = 32'h50413;
    ram[1755] = 32'h44052e23;
    ram[1756] = 32'h20000613;
    ram[1757] = 32'h593;
    ram[1758] = 32'h78513;
    ram[1759] = 32'h1c8000ef;
    ram[1760] = 32'h24a42a23;
    ram[1761] = 32'h46042023;
    ram[1762] = 32'h46042223;
    ram[1763] = 32'hc12083;
    ram[1764] = 32'h812403;
    ram[1765] = 32'h1010113;
    ram[1766] = 32'h8067;
    ram[1767] = 32'hff010113;
    ram[1768] = 32'h812423;
    ram[1769] = 32'h25452403;
    ram[1770] = 32'h912223;
    ram[1771] = 32'h112623;
    ram[1772] = 32'h50493;
    ram[1773] = 32'h41663;
    ram[1774] = 32'h100513;
    ram[1775] = 32'h240006f;
    ram[1776] = 32'h20442783;
    ram[1777] = 32'h79663;
    ram[1778] = 32'h20c42403;
    ram[1779] = 32'hfe9ff06f;
    ram[1780] = 32'h40593;
    ram[1781] = 32'h48513;
    ram[1782] = 32'he2dff0ef;
    ram[1783] = 32'hfe0516e3;
    ram[1784] = 32'hc12083;
    ram[1785] = 32'h812403;
    ram[1786] = 32'h412483;
    ram[1787] = 32'h1010113;
    ram[1788] = 32'h8067;
    ram[1789] = 32'hff010113;
    ram[1790] = 32'h812423;
    ram[1791] = 32'h1212023;
    ram[1792] = 32'h112623;
    ram[1793] = 32'h912223;
    ram[1794] = 32'h50913;
    ram[1795] = 32'h200413;
    ram[1796] = 32'h58463;
    ram[1797] = 32'h58413;
    ram[1798] = 32'h3092783;
    ram[1799] = 32'h745493;
    ram[1800] = 32'h79463;
    ram[1801] = 32'h845493;
    ram[1802] = 32'h1492583;
    ram[1803] = 32'h90513;
    ram[1804] = 32'hb485b3;
    ram[1805] = 32'he35ff0ef;
    ram[1806] = 32'hfff00793;
    ram[1807] = 32'h4050a63;
    ram[1808] = 32'h3092783;
    ram[1809] = 32'h20852703;
    ram[1810] = 32'h6079263;
    ram[1811] = 32'h849793;
    ram[1812] = 32'h40f407b3;
    ram[1813] = 32'h10437;
    ram[1814] = 32'hfff40413;
    ram[1815] = 32'h179793;
    ram[1816] = 32'h87f7b3;
    ram[1817] = 32'hf70433;
    ram[1818] = 32'h144783;
    ram[1819] = 32'h44503;
    ram[1820] = 32'hffff0737;
    ram[1821] = 32'h879793;
    ram[1822] = 32'ha787b3;
    ram[1823] = 32'h870713;
    ram[1824] = 32'he78733;
    ram[1825] = 32'h700693;
    ram[1826] = 32'he6e463;
    ram[1827] = 32'hfff00793;
    ram[1828] = 32'hc12083;
    ram[1829] = 32'h812403;
    ram[1830] = 32'h412483;
    ram[1831] = 32'h12903;
    ram[1832] = 32'h78513;
    ram[1833] = 32'h1010113;
    ram[1834] = 32'h8067;
    ram[1835] = 32'h749493;
    ram[1836] = 32'h40940433;
    ram[1837] = 32'h107b7;
    ram[1838] = 32'hfff78793;
    ram[1839] = 32'h241413;
    ram[1840] = 32'hf47433;
    ram[1841] = 32'h870433;
    ram[1842] = 32'h344783;
    ram[1843] = 32'h244503;
    ram[1844] = 32'hf0000737;
    ram[1845] = 32'h1879793;
    ram[1846] = 32'h1051513;
    ram[1847] = 32'ha787b3;
    ram[1848] = 32'h44503;
    ram[1849] = 32'ha787b3;
    ram[1850] = 32'h144503;
    ram[1851] = 32'h851513;
    ram[1852] = 32'ha787b3;
    ram[1853] = 32'h10000537;
    ram[1854] = 32'hfff50513;
    ram[1855] = 32'ha7f7b3;
    ram[1856] = 32'hf7dff06f;
    ram[1857] = 32'h50793;
    ram[1858] = 32'h7c703;
    ram[1859] = 32'h71663;
    ram[1860] = 32'h40a78533;
    ram[1861] = 32'h8067;
    ram[1862] = 32'h178793;
    ram[1863] = 32'hfedff06f;
    ram[1864] = 32'hc58633;
    ram[1865] = 32'h50793;
    ram[1866] = 32'hc59463;
    ram[1867] = 32'h8067;
    ram[1868] = 32'h5c703;
    ram[1869] = 32'h178793;
    ram[1870] = 32'h158593;
    ram[1871] = 32'hfee78fa3;
    ram[1872] = 32'hfe9ff06f;
    ram[1873] = 32'hc50633;
    ram[1874] = 32'h50793;
    ram[1875] = 32'hc79463;
    ram[1876] = 32'h8067;
    ram[1877] = 32'h178793;
    ram[1878] = 32'hfeb78fa3;
    ram[1879] = 32'hff1ff06f;
    ram[1880] = 32'h820017b7;
    ram[1881] = 32'h8ec7a703;
    ram[1882] = 32'h2071c63;
    ram[1883] = 32'hfff00513;
    ram[1884] = 32'h8067;
    ram[1885] = 32'h148493;
    ram[1886] = 32'h300e7;
    ram[1887] = 32'h4c503;
    ram[1888] = 32'h42303;
    ram[1889] = 32'hfe0518e3;
    ram[1890] = 32'h812403;
    ram[1891] = 32'hc12083;
    ram[1892] = 32'h412483;
    ram[1893] = 32'ha00513;
    ram[1894] = 32'h1010113;
    ram[1895] = 32'h30067;
    ram[1896] = 32'hff010113;
    ram[1897] = 32'h812423;
    ram[1898] = 32'h912223;
    ram[1899] = 32'h112623;
    ram[1900] = 32'h50493;
    ram[1901] = 32'h8ec78413;
    ram[1902] = 32'hfc5ff06f;
    ram[1903] = 32'h593;
    ram[1904] = 32'h92000537;
    ram[1905] = 32'h800006f;
    ram[1906] = 32'hff010113;
    ram[1907] = 32'h812423;
    ram[1908] = 32'h112623;
    ram[1909] = 32'h50413;
    ram[1910] = 32'h44503;
    ram[1911] = 32'h51a63;
    ram[1912] = 32'hc12083;
    ram[1913] = 32'h812403;
    ram[1914] = 32'h1010113;
    ram[1915] = 32'h8067;
    ram[1916] = 32'h140413;
    ram[1917] = 32'h64000ef;
    ram[1918] = 32'hfe1ff06f;
    ram[1919] = 32'hff010113;
    ram[1920] = 32'hfff00513;
    ram[1921] = 32'h112623;
    ram[1922] = 32'hb00fe0ef;
    ram[1923] = 32'hc00026f3;
    ram[1924] = 32'hc7b7;
    ram[1925] = 32'hb8078793;
    ram[1926] = 32'h2f6d6b3;
    ram[1927] = 32'hc0002773;
    ram[1928] = 32'h2f75733;
    ram[1929] = 32'h40d70733;
    ram[1930] = 32'hfea74ae3;
    ram[1931] = 32'h8067;
    ram[1932] = 32'hc0002573;
    ram[1933] = 32'hc7b7;
    ram[1934] = 32'hb8078793;
    ram[1935] = 32'h2f55533;
    ram[1936] = 32'h8067;
    ram[1937] = 32'h820017b7;
    ram[1938] = 32'h8ea7a823;
    ram[1939] = 32'h1300793;
    ram[1940] = 32'hf52623;
    ram[1941] = 32'h8067;
    ram[1942] = 32'h820017b7;
    ram[1943] = 32'h8f07a703;
    ram[1944] = 32'h872783;
    ram[1945] = 32'h87f793;
    ram[1946] = 32'hfe079ce3;
    ram[1947] = 32'ha72223;
    ram[1948] = 32'h513;
    ram[1949] = 32'h8067;
    ram[1950] = 32'h42204453;
    ram[1951] = 32'h6c746f6f;
    ram[1952] = 32'h6564616f;
    ram[1953] = 32'ha72;
    ram[1954] = 32'h6272;
    ram[1955] = 32'h6f6f622f;
    ram[1956] = 32'h69622e74;
    ram[1957] = 32'h6e;
    ram[1958] = 32'h2e2f2e2e;
    ram[1959] = 32'h72642f2e;
    ram[1960] = 32'h72657669;
    ram[1961] = 32'h64732f73;
    ram[1962] = 32'h5f64732f;
    ram[1963] = 32'h64726163;
    ram[1964] = 32'h632e;
    ram[1965] = 32'h61422221;
    ram[1966] = 32'h74732064;
    ram[1967] = 32'h22657461;
    ram[1968] = 32'h0;
    ram[1969] = 32'h45535341;
    ram[1970] = 32'h5452;
    ram[1971] = 32'h203a4453;
    ram[1972] = 32'h74696e49;
    ram[1973] = 32'h6d6f6320;
    ram[1974] = 32'h74656c70;
    ram[1975] = 32'h6465;
    ram[1976] = 32'h28282821;
    ram[1977] = 32'h746e6975;
    ram[1978] = 32'h745f3233;
    ram[1979] = 32'h72617429;
    ram[1980] = 32'h29746567;
    ram[1981] = 32'h33202620;
    ram[1982] = 32'h29;
    ram[1983] = 32'h0;
    ram[1984] = 32'h0;
    ram[1985] = 32'h0;
    ram[1986] = 32'h0;
    ram[1987] = 32'h0;
    ram[1988] = 32'h0;
    ram[1989] = 32'h0;
    ram[1990] = 32'h0;
end

// RAM write with byte enables
always @ (posedge clk_i)
begin
    if (ram_wr_w[0])
        ram[addr_w][7:0] <= ram_write_data_w[7:0];
    if (ram_wr_w[1])
        ram[addr_w][15:8] <= ram_write_data_w[15:8];
    if (ram_wr_w[2])
        ram[addr_w][23:16] <= ram_write_data_w[23:16];
    if (ram_wr_w[3])
        ram[addr_w][31:24] <= ram_write_data_w[31:24];

    ram_read_q <= ram[addr_w];
end

assign ram_read_data_w = ram_read_q;



endmodule
